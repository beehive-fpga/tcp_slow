module assembler_pipe (
     input clk
    ,input rst
);
endmodule   
